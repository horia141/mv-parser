module top;
   Data16to32 #(.Size(16))
   data ();
endmodule // top
